module LastConnect(
  input        clock,
  input        reset,
  input  [3:0] io_in,
  output [3:0] io_out
);
  assign io_out = 4'h4; // @[LastConnect.scala 14:10 LastConnect.scala 15:10 LastConnect.scala 16:10 LastConnect.scala 17:10]
endmodule
